`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.05.2022 22:14:11
// Design Name: 
// Module Name: fpm_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fpm_tb();
 reg [31:0]Num1,Num2;
 //wire [22:0]man_out;
 //wire [7:0]exp_out;
 //wire s_out;
 wire [31:0] final;
 
 fpm i1 (Num1,Num2,final);
 
 initial begin
 #0
 //3140000 and 26.43e-4
 Num1=32'b0_10010100_01111111010011010000000;
 Num2=32'b0_01110110_01011010011011000101110;
 //Sa=1'b0;Sb=1'b0;
 //Ea=8'b10010100; Eb=8'b01110110; 
 //Ma=23'b01111111010011010000000; Mb=23'b01011010011011000101110;
 #5
 //-2.78e-8 and 0.116e-11
 Num1=32'b1_01100101_11011101100110011011000;
 Num2=32'b0_01010111_01000110100000101100111;
 //Sa=1'b1; Sb=1'b0;
 //Ea=8'b01100101; Eb=8'b01010111;
// Ma=23'b11011101100110011011000; Mb=23'b01000110100000101100111;
#5
//-6.32e13 and -8.003e4
Num1=32'b1_10101100_11001011110101110010110;
Num2=32'b1_10001111_00111000100111100000000;

#5
Num1=32'b0_00000000_00000000000000000000000;
Num2=32'b01000000101000010000000000100000;

#5
// 4 and 5
Num1=32'b01000000100000000000000000000000;
Num2=32'b01000000101000000000000000000000;

#5$stop;


end
endmodule
